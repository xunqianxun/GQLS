module BTB (
    ports
);
    
endmodule